module tb;
  reg[7:0]din1,din2;
  reg[9:0]addr1,addr2;
  reg w_en1,w_en2;
  reg clk;
  wire [7:0]dout1,dout2;
  dual_ram_syn DUT(.*);
  initial begin
    clk=0;
    forever #5 clk=~clk;
  end
  initial begin
    clk=1;
    din1=8'd210;
    addr1=10'd1001;
    w_en1=1;
    din2=8'd210;
    addr2=10'd1010;
    w_en2=1;
    #10
    din1=8'd110;
    addr1=10'd999;
    w_en1=1;
    din2=8'd110;
    addr2=10'd888;
    w_en2=1;
   #10
    din1=8'd109;
    addr1=10'd777;
    w_en1=1;
    din2=8'd109;
    addr2=10'd666;
    w_en2=1;
   #10
    din1=8'd100;
    addr1=10'd999;
    w_en1=1;
    din2=8'd100;
    addr2=10'd698;
    w_en2=1;
   #10
    din1=8'd140;
    addr1=10'd1000;
    w_en1=1;
    din2=8'd140;
    addr2=10'd244;
    w_en2=1;
   #10
    din1=8'd178;
    addr1=10'd567;
    w_en1=1;
    din2=8'd178;
    addr2=10'd444;
    w_en2=1;
   #10
    din1=8'd220;
    addr1=10'd123;
    w_en1=1;
    din2=8'd220;
    addr2=10'd456;
    w_en2=1;
   #10
    din1=8'd250;
    addr1=10'd336;
    w_en1=1;
    din2=8'd250;
    addr2=10'd446;
    w_en2=1;
    #10
    din1=8'd210;
    addr1=10'd1001;
    w_en1=0;
    din2=8'd210;
    addr2=10'd1010;
    w_en2=0;
    #10
    din1=8'd110;
    addr1=10'd999;
    w_en1=0;
    din2=8'd110;
    addr2=10'd888;
    w_en2=0;
   #10
    din1=8'd109;
    addr1=10'd777;
    w_en1=0;
    din2=8'd109;
    addr2=10'd666;
    w_en2=0;
   #10
    din1=8'd100;
    addr1=10'd999;
    w_en1=0;
    din2=8'd100;
    addr2=10'd698;
    w_en2=0;
   #10
    din1=8'd140;
    addr1=10'd1000;
    w_en1=0;
    din2=8'd140;
    addr2=10'd244;
    w_en2=0;
   #10
    din1=8'd178;
    addr1=10'd567;
    w_en1=0;
    din2=8'd178;
    addr2=10'd444;
    w_en2=0;
   #10
    din1=8'd220;
    addr1=10'd123;
    w_en1=0;
    din2=8'd220;
    addr2=10'd456;
    w_en2=0;
   #10
    din1=8'd250;
    addr1=10'd336;
    w_en1=0;
    din2=8'd250;
    addr2=10'd446;
    w_en2=0;
    #10
    #600 $finish;
  end
    initial begin
      $monitor("time=%0t,INPUT VALUES:din1=%b,din2=%b,addr1=%b,addr2=%b,w_en1=%b,w_en2=%b,clk=%b, OUTPUT VALUES:dout1=%b,dout2=%b",$time,din1,din2,addr1,addr2,w_en1,w_en2,clk,dout1,dout2);
      $dumpfile("dual_ram_syn.vcd");
      $dumpvars;
      end
endmodule
